module neural_network_top (
    input CLOCK_50,
    input [1:0] KEY,   // Start signal (active low)
    input [9:0] SW,
	 input i_RX_Serial,
    output [9:0] LEDR, // LEDs for state indication
    output [6:0] HEX0  // 7-segment display for output
);

    // Internal signals
    wire clk;
    wire clk_slow;
    wire start;
    wire resetn;
    wire done;
    wire [3:0] argmax_output;
	 wire [31:0] mm1_debug_data;
	 wire [31:0] mm2_debug_data;
	 wire [31:0] mm4_debug_data;
	 wire [31:0] matrix1_data;
    
    // State signals
    wire [3:0] current_state;
    wire [3:0] next_state;
    
    // Clock divider instance
    clock_divider clk_div (
        .clk_in(CLOCK_50),
        .clk_out(clk_slow),
        .DIVISOR(32'd500)  // Adjust this value to change clock speed
    );

    // Assign clock, start and reset
    assign clk = clk_slow;  // Use the slower clock
    assign start = ~KEY[0]; // KEY[0] is used for start
    assign resetn = SW[0];

    assign LEDR[9] = start;  // Shows if start is active
    assign LEDR[3:0] = current_state;  // Shows current state in binary

    // Neural network instance
    neural_network nn (
        .clk(clk),
        .resetn(resetn),
        .start(start),
        .rx_serial(i_RX_Serial),
        .done(done),
        .current_state(current_state),
        .next_state(next_state),
        .argmax_output(argmax_output)
    );
 
	 
	 DisplayNum display_hex(
		  .num(argmax_output),
		  .hex(HEX0)
	 );
	 
	 image_memory weight_mem1(
        .address(5),
        .data_out(matrix1_data)
    );

endmodule
